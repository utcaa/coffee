Email|First Name|Last Name|Preferred Name|School|Grad year|Majors|Years of Wokring Experience|Employers|current role|current industry|current function
Jennifer.zhu@tdam.com|Jennifer|Zhu||UofT|2010|Finance|>5 years|TD Asset Management|Associate|Investment Management|Investment Management
jordanhwh@gmail.com|Steven|He||UofT|2016|Engineering Science|1-3 years|Point72, RBC Capital Markets|Associate|Investment Management|Investment Management
herrydai.hd@gmail.com|Herry|Dai||UofT|2012|Finance|More than 5 years|Canada Post Pension, OBSI, Citigroup, Garrison Hill|Manager/Supervisor|Investment Management|Investment Management
sihang.lin@gmail.com|Leo|Lin||UofT|2011|B.Com, accounting specialist|More than 5 years|Osisko Mining, Largardere, Corsa Coal, EY|Manager/Supervisor|Exact Minerals/Metals|Accounting
ziqing.mt@gmail.com|Ziqing|Tang|Michael|UofT|2013|EngSci|1-3 years|Waratah|Analyst|Investment Management|Investment Management
seanroylv@hotmail.com|Cheng|Lu||UofT|2013|Finance and Economics|3-5 years|National Bank of Canada, Canaccord Genuity, OBSI|Analyst|Investment Banking/Brokerage/Securities|Investment Banking
hepy1227@hotmail.com|Peiyang|He||UofT|2014|statistics |3-5 years|Amazon, TD Bank, RSA Canada|Analyst, Data scientist|Retail|Product Management, Data Science
haosheng.li@hotmail.com|Haosheng|Li||New York University - Courant Institute of Mathematical Sciences|2016|Mathematics in Finance|1-3 years|Alignvest Investment Management, Morneau Shepell, PwC Canada|Analyst|Investment Management|Investment Management
Jackson.mei@td.com|Jackson|Mei||UofT|2012|Management|More than 5 years|TD, BCE, AGF|Manager/Supervisor|Diversified Financial Services|Finance
Zhenyu.luo@mail.utoronto.ca|Dennis|Luo||UofT|2016|Mathematical Finance|1-3 years|University of Toronto Asset Management|Analyst|Investment Management|Investment Management
bei.liu.utsc@gmail.com|Cindy |Liu||UofT|2017|Master of Mangement and Professional Accounting|1-3 years|Fuller Landau LLP (current), Manulife, TD, Ontario Ministry of Finance|Analyst|Accounting|Accounting
mabelmwang@gmail.com|Mable|Wang||UofT|2012|Commerce|> 5 years|Bank of Nova Scotia|Manager/Supervior|Transportation Services|Finance - Group Treasury
chixiao429429@hotmail.com|Shawn|Xiao||UofT|2011|Engineering|> 5 years|ASC EBS|Director/VP|Entertainment/Leisure|General Management
Michelle.duan19@rotman.utoronto.ca|Michelle|Duan||University of Calgary|2012|Chemical Engineering|>5 years|Rotman MBA, Trans Canada|MBA candidate|Education|Engineering
cindy.xu0112@gmail.com|Yunying|Xu|Cindy|UofT|2016|Accounting|1-3 years|Accountable Solutions|Junior Accountant|Accounting|Accounting
John.hanfeng@gmail.com|John|Guo||UofT|2016|Mechanical Engineering|1-3 years|Acculogic Inc. (current), Shadefx Canopies Inc., CardioMed Supplies Inc.|Associate|Manufacturing|Engineering
sylvialiu2012@gmail.com|Xi|Liu|Sylvia|McMaster University|2015|Finance|1-3 years|CDLSI, H&R Block|Analyst|Auto|Service Marketing, Car Lease
amychen.education@gmail.com|Amy|Chen||UofT|2017|Political Science and History|1-3 years|Top Hat, University of Toronto, Sensors Quality Management Inc.|Associate, Postgraduate Journalism student|Media, Journalism|Nonprofit, Journalist
Jerryfeng2@gmail.com|Jerry|Feng||UofT|2016|Master of Financial Economics|1-3 years|Deloitte, TD Bank Group, University of Toronto Asset Management Corp.|Associate|Risk Management|Finance
yizhi_zhang@icloud.com|yizhi|zhang|university of ottawa|UofT|2015|system science|3-5 years|eq works, university of ottawa|Associate, designer|Software, designer|Strategic Planning, Designer and developer
mobyrobin@gmail.com|Yanlin|Sun|Moby|UofT|2012|Management & Accounting|More than 5 years|Shaw Communications|Analyst|Telecom|Accounting
alice.h.luo@gmail.com|Alice|Luo||U of T (Rotman MBA)|2017|Strategy|1-3 years|"Self-employed, boutique mgmt consulting firm
, EY, UBS"|Associate|Consulting|Consulting
kwokwil0323@gmail.com|William|Kwok||UofT|2014|Industrial engineering|3-5 years|EY, Accenture, Scotiabank|Associate|Consulting|Consulting
Yohancong@gmail.com|Yohan|Cong||UofT|2013|Accounting|3-5 years|EY, MNP, Auditor General of Canada|Manager/Supervisor|Accounting|Accounting
christyz0406@gmail.com|Christy|Zhang||UofT|2015|Accounting|1-3 years|Accountable Solutions Accounting Professional Corporation|Manager/Supervisor|Accounting|Accounting
Yizhu.wang@mail.utoronto.ca|Janet|Wang||UofT Scarborough|2012|Management and Human Resources|More than 5 years|Sun Life Financial, Rogers Communications Inc|Associate|Insurance|Human Resources
Kx3@ntrs.com|Kiana|Xu||UofT, Rotman Commerce|2012|Finance and Economics|More than 5 years|Northern Trust Asset Management, BNY Mellon Wealth Management|Analyst|Investment Management|Investment Management
arielw22@hotmail.com|Ariel|Wang||UofT|2015|statistics and Economics|1-3 years|RBC Capital Markets|Analyst|Risk Management|Finance, Data Management
pete.wong@utoronto.ca|Peter|Wong||UofT|2004|Genetics/Economics|More than 5 years|University of Toronto|Associate, Senior Auditor|Education|Accounting
alexyucanada@gmail.com|思谦|余||Georgian College|2016|Computer Science|1-3 years|UPS|Associate|Transportation Services|Business Development
evangelinkoko1482@Hotmail.com|Evangeline|Zhou||UofT|2012|Management and Humanities|3-5 years|Toronto Mandarin School|Analyst|Education|Administration
Sallylyq0126@gmail.com|Sally|Li||UofT|2015|Political Science Specialist|1-3 years|Golden Voice English|Analyst, Coordinator|Data Analytics|Operations
james.zefang.li@gmail.com|James|Li||UofT|2015|Materials Engineering|1-3 years|Shawcor|Associate|Energy|Engineering
lhy_james@hotmail.com|Haoyang|Liang||U of T|2012|csc & sta|More than 5 years|DBRS, Oracle, Amazon, Wherego|C-Level (CEO, CFO, COO, etc)|Computer - Related Services|General Management
loewe.ke@kesolutions.ca|Loewe|Ke||University of Waterloo|2011|Actuarial Science and Computer Science|More than 5 years|KE Solutions|C-Level (CEO, CFO, COO, etc)|Data Analytics|Consulting
jyang.xia@gmail.com|Jake|Xia||Uoft and ryerson|2011|Dietitian and food science/nutritional science|More than 5 years|Candian food Inspection agency|Associate/Analyst|Government|Auditing
