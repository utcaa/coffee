UTmail|First Name|Last Name|Preferred Name|School|Grad (expected) year|Majors|Where have you worked|Recent/Interested Role|Recent/Interested Industry|Interests&Career Plan|Challenges|Coffe chat goals| want to be paired up with|preferred location|# of chat avaiability|additional comments||Professional Matching|potential match|Responsibile|Notes|professional list|Dates Added
janet.tan@mail.utoronto.ca|simin|tan|janet|U of T|2018|public accounting|Geodis supply chain|Accounting|Accounting|I am going to study in the master of taxation program at the University of Waterloo and I planning to acquire an accounting related position in the future|Building a resume,Looking for a job|1. build network 2. ask for career advice 3.find job opportunities|accounting professional|downtown|1|||sihang.lin@gmail.com|||||May 2018
Michelle.duan19@rotman.utoronto.ca|Michelle|Duan||U of T|2019|Rotman MBA|Trans Canada, Johnson & Johnson|Consulting|Health Services|Interested in healthcare consulting and strategy|Looking for a mentor|1. mentorship 2. industry development|any industry|downtown|5|||unmatched||Alice will follow up|||May 2018
jiajie.li19@rotman.utoronto.ca|jiajie|Li|Jack|U of T|2019|Rotman MBA|Nestle|Entrepreneurship|TMT|Entrepreneurship. Build a startup in China|Looking for a mentor|1.looking for mentors 2. Looking for technical people 3. build network|Technology, founder of startup if possible|downtown|1-2|I would appreciate it if you could tell me how you match us||unmatched||Alice will follow up|done|alice.h.luo@gmail.com|May 2018
naiying.zhu@mail.utoronto.ca|Naiying|Zhu||U of T|2019|Economics and Statistics||Investment Banking|Investment Banking/Brokerage/Securities|Consulting and Investment Bank|1. build a resume 2.looking for a job 3.network with others|1.build network 2.Ask for career advice|Banking, Consulting|downtown|5|||jordanhwh@gmail.com|||||May 2018
juntian.li@mail.utoronto.ca|Juntian|Li||U of T|2019|Master of Global Affairs|Ministry of Economic Growth and Development|Busnisess Develpoment|Government|Management and Innovation.|1. build a resume 2.looking for a mentor 3. looking for a job 3.studying 4. studying|1. build network 2.find job opportunities 3. ask for career advice|N/A|DT, Mississauga|1|||alice.h.luo@gmail.com|||||May 2018
jingrui.gu@mail.utoronto.ca|Serena(Jingrui)|Gu|Serena|UTSC|2021|Mental Health Studies||Human Resources|Psychology, Human Resources|1. Mental Health 2. psychologist\psychiatrist 3. HR|1. Looking for a mentor 2. Looking for a job 3. Career expectation and choices|1. build networks 2.ask for career advice 3. ask about the future of fields inluding psychology and HR|professions in psychology or HR or seniors student in these fields|Scarborough��Downtown|many|||Yizhu.wang@mail.utoronto.ca|||||May 2018
boey.li@mail.utoronto.ca|Boey|Li||U of T|2020|Rotman Commerce Public Accounting||Accounting|Accounting|N/A|N/A|N/A|N/A|N/A|N/A|||christyz0406@gmail.com|||||May 2018
yuning.zhang@mail.utoronto.ca|Yuning|Zhang|Jessica|U of T|2018|Rotman Commerce- Finance& Economy|IBM, U of T, Bluekey Education|Operations|Diversifieed Financial Services|Interests: Finance, Tecnology, Non-Profit (Marketing), Consulting Career Plan: full time roles related to Finance & Technology, part-time/volunteer in non-profit => UN oversea volunteering => MBA => consulting or Non-profit|1. build a resume 2. Looking for a mentor 3. Looking for a job|1. Ask for career advice 2. Find job opportunities 3. Build network|Fin Tech|Downtown, North York, Markham|As many as possible|||herrydai.hd@gmail.com|||||May 2018
Christina.guo@mail.utoronto.ca|Christina|Guo|Clover|U of T|2017|Statistic|CIBC|Finance|Analyst|Business analyst|1. looking for a mentor 2. looking for a job|1.Ask for career advice 2. Build networking 3. Find job|Banker|North York|2-3|||Kx3@ntrs.com|||||May 2018
huanyu.jiang@mail.utoronto.ca|mya|jiang|uoft|2021|engineering|New oriental education inc|Energy|Enineering|Be an engineer |Building a resume, Looking for a mentor, Looking for a job|Build network and get advice|Professionals in engineering, biomedical, aerospace and finance|A month|A month|A month|Downtown|||||||May 2018
