student_id|interest_industry_id|interest_role_id|goal|comments|challenge|location_id
c99752c5-9a57-417e-8c61-d4e031f8680f|9|1|go test2|cm test2|ch test2|4089
9ed2d02f-b77d-4b0c-bc4b-243d83b19c97|1|1|go test1|cm test1|ch test1|4089