student_id|interest_industry_id|interest_role_id|goal|comments|challenge|location_id
1|1|1|go test1|cm test1|ch test1|4089
1|1|1|go test2|cm test2|ch test2|4089